package core_eei;
    localparam int unsigned MEM_DATA_WIDTH = 32;
endpackage
