

module core_top
    import core_eei::*;
;
    core___membus_if__eei_MEM_DATA_WIDTH__20 membus ();
endmodule
